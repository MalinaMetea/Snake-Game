module characters_ROM
   (
    input wire clk_25,
    input wire [10:0] address,
    output reg [7:0] data
   );
   
reg [10:0] address_reg; 

always @(posedge clk_25) 
begin
    address_reg <= address;
end
	  
always @(*)
begin
    case (address_reg) // daca folosesc direct addr nu arata clar textul)  	  
             11'h000: data = 8'b00000000; // 
             11'h001: data = 8'b00000000; // 
             11'h002: data = 8'b00000000; // 
             11'h003: data = 8'b00000000; // 
             11'h004: data = 8'b00000000; // 
             11'h005: data = 8'b00000000; // 
             11'h006: data = 8'b00000000; // 
             11'h007: data = 8'b00000000; // 
             11'h008: data = 8'b00000000; // 
             11'h009: data = 8'b00000000; // 
             11'h00a: data = 8'b00000000; // 
             11'h00b: data = 8'b00000000; // 
             11'h00c: data = 8'b00000000; // 
             11'h00d: data = 8'b00000000; // 
             11'h00e: data = 8'b00000000; // 
             11'h00f: data = 8'b00000000; // 
             
    //code x01
             11'h010: data = 8'b00000000; // 
             11'h011: data = 8'b00000000; // 
             11'h012: data = 8'b01111100; //  *****
             11'h013: data = 8'b11000110; // **   **
             11'h014: data = 8'b11000110; // **   **
             11'h015: data = 8'b11001110; // **  ***
             11'h016: data = 8'b11011110; // ** ****
             11'h017: data = 8'b11110110; // **** **
             11'h018: data = 8'b11100110; // ***  **
             11'h019: data = 8'b11000110; // **   **
             11'h01a: data = 8'b11000110; // **   **
             11'h01b: data = 8'b01111100; //  *****
             11'h01c: data = 8'b00000000; // 
             11'h01d: data = 8'b00000000; // 
             11'h01e: data = 8'b00000000; // 
             11'h01f: data = 8'b00000000; // 
             
    //code x02
             11'h020: data = 8'b00000000; // 
             11'h021: data = 8'b00000000; // 
             11'h022: data = 8'b00011000; // 
             11'h023: data = 8'b00011100; // 
             11'h024: data = 8'b00011110; //    **
             11'h025: data = 8'b00011000; //   ***
             11'h026: data = 8'b00011000; //  ****
             11'h027: data = 8'b00011000; //    **
             11'h028: data = 8'b00011000; //    **
             11'h029: data = 8'b00011000; //    **
             11'h02a: data = 8'b00011000; //    **
             11'h02b: data = 8'b01111110; //    **
             11'h02c: data = 8'b00000000; //    **
             11'h02d: data = 8'b00000000; //  ******
             11'h02e: data = 8'b00000000; // 
             11'h02f: data = 8'b00000000; // 
             
    //code x03
             11'h030: data = 8'b00000000; // 
             11'h031: data = 8'b00000000; // 
             11'h032: data = 8'b00111110; //  *****
             11'h033: data = 8'b01100011; // **   **
             11'h034: data = 8'b01100000; //      **
             11'h035: data = 8'b00110000; //     **
             11'h036: data = 8'b00011000; //    **
             11'h037: data = 8'b00001100; //   **
             11'h038: data = 8'b00000110; //  **
             11'h039: data = 8'b00000011; // **
             11'h03a: data = 8'b01100011; // **   **
             11'h03b: data = 8'b01111111; // *******
             11'h03c: data = 8'b00000000; // 
             11'h03d: data = 8'b00000000; // 
             11'h03e: data = 8'b00000000; // 
             11'h03f: data = 8'b00000000; // 
             
    //code x04
             11'h040: data = 8'b00000000; // 
             11'h041: data = 8'b00000000; // 
             11'h042: data = 8'b00111110; //  *****
             11'h043: data = 8'b01100011; // **   **
             11'h044: data = 8'b01100000; //      **
             11'h045: data = 8'b01100000; //      **
             11'h046: data = 8'b00111100; //   ****
             11'h047: data = 8'b01100000; //      **
             11'h048: data = 8'b01100000; //      **
             11'h049: data = 8'b01100000; //      **
             11'h04a: data = 8'b01100011; // **   **
             11'h04b: data = 8'b00111110; //  *****
             11'h04c: data = 8'b00000000; // 
             11'h04d: data = 8'b00000000; // 
             11'h04e: data = 8'b00000000; // 
             11'h04f: data = 8'b00000000; // 
             
    //code x05
             11'h050: data = 8'b00000000; // 
             11'h051: data = 8'b00000000; // 
             11'h052: data = 8'b00110000; //     **
             11'h053: data = 8'b00111000; //    ***
             11'h054: data = 8'b00111100; //   ****
             11'h055: data = 8'b00110110; //  ** **
             11'h056: data = 8'b00110011; // **  **
             11'h057: data = 8'b01111111; // *******
             11'h058: data = 8'b00110000; //     **
             11'h059: data = 8'b00110000; //     **
             11'h05a: data = 8'b00110000; //     **
             11'h05b: data = 8'b01111000; //    ****
             11'h05c: data = 8'b00000000; // 
             11'h05d: data = 8'b00000000; // 
             11'h05e: data = 8'b00000000; // 
             11'h05f: data = 8'b00000000; // 
    
    //code x06
             11'h060: data = 8'b00000000; // 
             11'h061: data = 8'b00000000; // 
             11'h062: data = 8'b01111111; // *******
             11'h063: data = 8'b00000011; // **
             11'h064: data = 8'b00000011; // **
             11'h065: data = 8'b00000011; // **
             11'h066: data = 8'b00111111; // ******
             11'h067: data = 8'b01100000; //      **
             11'h068: data = 8'b01100000; //      **
             11'h069: data = 8'b01100000; //      **
             11'h06a: data = 8'b01100011; // **   **
             11'h06b: data = 8'b00111110; //  *****
             11'h06c: data = 8'b00000000; // 
             11'h06d: data = 8'b00000000; // 
             11'h06e: data = 8'b00000000; // 
             11'h06f: data = 8'b00000000; // 
    
    //code x07
             11'h070: data = 8'b00000000; // 
             11'h071: data = 8'b00000000; // 
             11'h072: data = 8'b00011100; //   ***
             11'h073: data = 8'b00000110; //  **
             11'h074: data = 8'b00000011; // **
             11'h075: data = 8'b00000011; // **
             11'h076: data = 8'b00111111; // ******
             11'h077: data = 8'b01100011; // **   **
             11'h078: data = 8'b01100011; // **   **
             11'h079: data = 8'b01100011; // **   **
             11'h07a: data = 8'b01100011; // **   **
             11'h07b: data = 8'b00111110; //  *****
             11'h07c: data = 8'b00000000; // 
             11'h07d: data = 8'b00000000; // 
             11'h07e: data = 8'b00000000; // 
             11'h07f: data = 8'b00000000; // 
    
    //code x08
             11'h080: data = 8'b00000000; // 
             11'h081: data = 8'b00000000; // 
             11'h082: data = 8'b01111111; // *******
             11'h083: data = 8'b01100000; // **   **
             11'h084: data = 8'b01100000; //      **
             11'h085: data = 8'b01100000; //      **
             11'h086: data = 8'b00110000; //     **
             11'h087: data = 8'b00011000; //    **
             11'h088: data = 8'b00001100; //   **
             11'h089: data = 8'b00001100; //   **
             11'h08a: data = 8'b00001100; //   **
             11'h08b: data = 8'b00001100; //   **
             11'h08c: data = 8'b00000000; // 
             11'h08d: data = 8'b00000000; // 
             11'h08e: data = 8'b00000000; // 
    
    //code x09
             11'h090: data = 8'b00000000; // 
             11'h091: data = 8'b00000000; // 
             11'h092: data = 8'b01111100; //  *****
             11'h093: data = 8'b11000110; // **   **
             11'h094: data = 8'b11000110; // **   **
             11'h095: data = 8'b11000110; // **   **
             11'h096: data = 8'b01111100; //  *****
             11'h097: data = 8'b11000110; // **   **
             11'h098: data = 8'b11000110; // **   **
             11'h099: data = 8'b11000110; // **   **
             11'h09a: data = 8'b11000110; // **   **
             11'h09b: data = 8'b01111100; //  *****
             11'h09c: data = 8'b00000000; // 
             11'h09d: data = 8'b00000000; // 
             11'h09e: data = 8'b00000000; // 
             11'h09f: data = 8'b00000000; // 
    
    //code x0a
             11'h0a0: data = 8'b00000000; // 
             11'h0a1: data = 8'b00000000; // 
             11'h0a2: data = 8'b00111110; //  *****
             11'h0a3: data = 8'b01100011; // **   **
             11'h0a4: data = 8'b01100011; // **   **
             11'h0a5: data = 8'b01100011; // **   **
             11'h0a6: data = 8'b01111110; //  ******
             11'h0a7: data = 8'b01100000; //      **
             11'h0a8: data = 8'b01100000; //      **
             11'h0a9: data = 8'b01100000; //      **
             11'h0aa: data = 8'b00110000; //     **
             11'h0ab: data = 8'b00011110; //  ****
             11'h0ac: data = 8'b00000000; // 
             11'h0ad: data = 8'b00000000; // 
             11'h0ae: data = 8'b00000000; // 
             11'h0af: data = 8'b00000000; // 		 
    
    //code x0b
             11'h0b0: data = 8'b00000000; // 
             11'h0b1: data = 8'b00000000; // 
             11'h0b2: data = 8'b00010000; //    *
             11'h0b3: data = 8'b00111000; //   ***
             11'h0b4: data = 8'b01101100; //  ** **
             11'h0b5: data = 8'b11000110; // **   **
             11'h0b6: data = 8'b11000110; // **   **
             11'h0b7: data = 8'b11111110; // *******
             11'h0b8: data = 8'b11000110; // **   **
             11'h0b9: data = 8'b11000110; // **   **
             11'h0ba: data = 8'b11000110; // **   **
             11'h0bb: data = 8'b11000110; // **   **
             11'h0bc: data = 8'b00000000; // 
             11'h0bd: data = 8'b00000000; // 
             11'h0be: data = 8'b00000000; // 
             11'h0bf: data = 8'b00000000; // 
    
    //code x0c
             11'h0c0: data = 8'b00000000; // 
             11'h0c1: data = 8'b00000000; // 
             11'h0c2: data = 8'b11111100; // ******
             11'h0c3: data = 8'b01100110; //  **  **
             11'h0c4: data = 8'b01100110; //  **  **
             11'h0c5: data = 8'b01100110; //  **  **
             11'h0c6: data = 8'b01111100; //  *****
             11'h0c7: data = 8'b01100110; //  **  **
             11'h0c8: data = 8'b01100110; //  **  **
             11'h0c9: data = 8'b01100110; //  **  **
             11'h0ca: data = 8'b01100110; //  **  **
             11'h0cb: data = 8'b11111100; // ******
             11'h0cc: data = 8'b00000000; // 
             11'h0cd: data = 8'b00000000; // 
             11'h0ce: data = 8'b00000000; // 
             11'h0cf: data = 8'b00000000; // 
             
    //code x0d
             11'h0d0: data = 8'b00000000; // 
             11'h0d1: data = 8'b00000000; // 
             11'h0d2: data = 8'b00111100; //   ****
             11'h0d3: data = 8'b01100110; //  **  **
             11'h0d4: data = 8'b01000011; // **    *
             11'h0d5: data = 8'b00000011; // **
             11'h0d6: data = 8'b00000011; // **
             11'h0d7: data = 8'b00000011; // **
             11'h0d8: data = 8'b00000011; // **
             11'h0d9: data = 8'b01000011; // **    *
             11'h0da: data = 8'b01100110; //  **  **
             11'h0db: data = 8'b01111110; //   ****
             11'h0dc: data = 8'b00000000; // 
             11'h0dd: data = 8'b00000000; // 
             11'h0de: data = 8'b00000000; // 
             11'h0df: data = 8'b00000000; // 
    
    //code x0e 
             11'h0e0: data = 8'b00000000; // 
             11'h0e1: data = 8'b00000000; // 
             11'h0e2: data = 8'b11111000; // *****
             11'h0e3: data = 8'b01101100; //  ** **
             11'h40e: data = 8'b01100110; //  **  **
             11'h0e5: data = 8'b01100110; //  **  **
             11'h0e6: data = 8'b01100110; //  **  **
             11'h0e7: data = 8'b01100110; //  **  **
             11'h0e8: data = 8'b01100110; //  **  **
             11'h0e9: data = 8'b01100110; //  **  **
             11'h0ea: data = 8'b01101100; //  ** **
             11'h0eb: data = 8'b11111000; // *****
             11'h0ec: data = 8'b00000000; // 
             11'h0ed: data = 8'b00000000; // 
             11'h0ee: data = 8'b00000000; // 
             11'h0ef: data = 8'b00000000; // 
    
    //code x0f
             11'h0f0: data = 8'b00000000; // 
             11'h0f1: data = 8'b00000000; // 
             11'h0f2: data = 8'b01111111; // *******
             11'h0f3: data = 8'b01100110; //  **  **
             11'h0f4: data = 8'b01000110; //  **   *
             11'h0f5: data = 8'b00010110; //  ** *
             11'h0f6: data = 8'b00011110; //  ****
             11'h0f7: data = 8'b00010110; //  ** *
             11'h0f8: data = 8'b00000110; //  **
             11'h0f9: data = 8'b01000110; //  **   *
             11'h0fa: data = 8'b01100110; //  **  **
             11'h0fb: data = 8'b01111111; // *******
             11'h0fc: data = 8'b00000000; // 
             11'h0fd: data = 8'b00000000; // 
             11'h0fe: data = 8'b00000000; // 
             11'h0ff: data = 8'b00000000; // 
    
    //code x10
             11'h100: data = 8'b00000000; // 
             11'h101: data = 8'b00000000; // 
             11'h102: data = 8'b11111110; // *******
             11'h103: data = 8'b01100110; //  **  **
             11'h104: data = 8'b01100010; //  **   *
             11'h105: data = 8'b01101000; //  ** *
             11'h106: data = 8'b01111000; //  ****
             11'h107: data = 8'b01101000; //  ** *
             11'h108: data = 8'b01100000; //  **
             11'h109: data = 8'b01100000; //  **
             11'h10a: data = 8'b01100000; //  **
             11'h10b: data = 8'b11110000; // ****
             11'h10c: data = 8'b00000000; // 
             11'h10d: data = 8'b00000000; // 
             11'h10e: data = 8'b00000000; // 
             11'h10f: data = 8'b00000000; // 
    
    //code x11
             11'h110: data = 8'b00000000; // 
             11'h111: data = 8'b00000000; // 
             11'h112: data = 8'b00111100; //   ****
             11'h113: data = 8'b01100110; //  **  **
             11'h114: data = 8'b01000011; // **    *
             11'h115: data = 8'b00000011; // **
             11'h116: data = 8'b00000011; // **
             11'h117: data = 8'b01111011; // ** ****
             11'h118: data = 8'b01100011; // **   **
             11'h119: data = 8'b01100011; // **   **
             11'h11a: data = 8'b01100110; //  **  **
             11'h11b: data = 8'b01011100; //   *** *
             11'h11c: data = 8'b00000000; // 
             11'h11d: data = 8'b00000000; // 
             11'h11e: data = 8'b00000000; // 
             11'h11f: data = 8'b00000000; // 
             
    //code x12
             11'h120: data = 8'b00000000; // 
             11'h121: data = 8'b00000000; // 
             11'h122: data = 8'b11000110; // **   **
             11'h123: data = 8'b11000110; // **   **
             11'h124: data = 8'b11000110; // **   **
             11'h125: data = 8'b11000110; // **   **
             11'h126: data = 8'b11111110; // *******
             11'h127: data = 8'b11000110; // **   **
             11'h128: data = 8'b11000110; // **   **
             11'h129: data = 8'b11000110; // **   **
             11'h12a: data = 8'b11000110; // **   **
             11'h12b: data = 8'b11000110; // **   **
             11'h12c: data = 8'b00000000; // 
             11'h12d: data = 8'b00000000; // 
             11'h12e: data = 8'b00000000; // 
             11'h12f: data = 8'b00000000; // 
    
    //code x13
             11'h130: data = 8'b00000000; // 
             11'h131: data = 8'b00000000; // 
             11'h132: data = 8'b00111100; //   ****
             11'h133: data = 8'b00011000; //    **
             11'h134: data = 8'b00011000; //    **
             11'h135: data = 8'b00011000; //    **
             11'h136: data = 8'b00011000; //    **
             11'h137: data = 8'b00011000; //    **
             11'h138: data = 8'b00011000; //    **
             11'h139: data = 8'b00011000; //    **
             11'h13a: data = 8'b00011000; //    **
             11'h13b: data = 8'b00111100; //   ****
             11'h13c: data = 8'b00000000; // 
             11'h13d: data = 8'b00000000; // 
             11'h13e: data = 8'b00000000; // 
             11'h13f: data = 8'b00000000; // 
    
    //code x14 
             11'h140: data = 8'b00000000; // 
             11'h141: data = 8'b00000000; // 
             11'h142: data = 8'b00011110; //    ****
             11'h143: data = 8'b00001100; //     **
             11'h144: data = 8'b00001100; //     **
             11'h145: data = 8'b00001100; //     **
             11'h146: data = 8'b00001100; //     **
             11'h147: data = 8'b00001100; //     **
             11'h148: data = 8'b11001100; // **  **
             11'h149: data = 8'b11001100; // **  **
             11'h14a: data = 8'b11001100; // **  **
             11'h14b: data = 8'b01111000; //  ****
             11'h14c: data = 8'b00000000; // 
             11'h14d: data = 8'b00000000; // 
             11'h14e: data = 8'b00000000; // 
             11'h14f: data = 8'b00000000; // 
    
    //code x15  
             11'h150: data = 8'b00000000; // 
             11'h151: data = 8'b00000000; // 
             11'h152: data = 8'b11100110; // ***  **
             11'h153: data = 8'b01100110; //  **  **
             11'h154: data = 8'b01100110; //  **  **
             11'h155: data = 8'b01101100; //  ** **
             11'h156: data = 8'b01111000; //  ****
             11'h157: data = 8'b01111000; //  ****
             11'h158: data = 8'b01101100; //  ** **
             11'h159: data = 8'b01100110; //  **  **
             11'h15a: data = 8'b01100110; //  **  **
             11'h15b: data = 8'b11100110; // ***  **
             11'h15c: data = 8'b00000000; // 
             11'h15d: data = 8'b00000000; // 
             11'h15e: data = 8'b00000000; // 
             11'h15f: data = 8'b00000000; // 
    
    //code x16 
             11'h160: data = 8'b00000000; // 
             11'h161: data = 8'b00000000; // 
             11'h162: data = 8'b00001111; // ****
             11'h163: data = 8'b00000110; //  **
             11'h164: data = 8'b00000110; //  **
             11'h165: data = 8'b00000110; //  **
             11'h166: data = 8'b00000110; //  **
             11'h167: data = 8'b00000110; //  **
             11'h168: data = 8'b00000110; //  **
             11'h169: data = 8'b01000110; //  **   *
             11'h16a: data = 8'b01100110; //  **  **
             11'h16b: data = 8'b01111111; // *******
             11'h16c: data = 8'b00000000; // 
             11'h16d: data = 8'b00000000; // 
             11'h16e: data = 8'b00000000; // 
             11'h16f: data = 8'b00000000; // 
    
    //code x17  
             11'h170: data = 8'b00000000; // 
             11'h171: data = 8'b00000000; // 
             11'h172: data = 8'b11000011; // **    **
             11'h173: data = 8'b11100111; // ***  ***
             11'h174: data = 8'b11111111; // ********
             11'h175: data = 8'b11111111; // ********
             11'h176: data = 8'b11011011; // ** ** **
             11'h177: data = 8'b11000011; // **    **
             11'h178: data = 8'b11000011; // **    **
             11'h179: data = 8'b11000011; // **    **
             11'h17a: data = 8'b11000011; // **    **
             11'h17b: data = 8'b11000011; // **    **
             11'h17c: data = 8'b00000000; // 
             11'h17d: data = 8'b00000000; // 
             11'h17e: data = 8'b00000000; // 
             11'h17f: data = 8'b00000000; // 
    
    //code x18
             11'h180: data = 8'b00000000; // 
             11'h181: data = 8'b00000000; // 
             11'h182: data = 8'b01100011; // **   **
             11'h183: data = 8'b01100111; // ***  **
             11'h184: data = 8'b01101111; // **** **
             11'h185: data = 8'b01111111; // *******
             11'h186: data = 8'b01110111; // ** ****
             11'h187: data = 8'b01100111; // **  ***
             11'h188: data = 8'b01100011; // **   **
             11'h189: data = 8'b01100011; // **   **
             11'h18a: data = 8'b01100011; // **   **
             11'h18b: data = 8'b01100011; // **   **
             11'h18c: data = 8'b00000000; // 
             11'h18d: data = 8'b00000000; // 
             11'h18e: data = 8'b00000000; // 
             11'h18f: data = 8'b00000000; // 
    
    //code x19 
             11'h190: data = 8'b00000000; // 
             11'h191: data = 8'b00000000; // 
             11'h192: data = 8'b01111100; //  *****
             11'h193: data = 8'b11000110; // **   **
             11'h194: data = 8'b11000110; // **   **
             11'h195: data = 8'b11000110; // **   **
             11'h196: data = 8'b11000110; // **   **
             11'h197: data = 8'b11000110; // **   **
             11'h198: data = 8'b11000110; // **   **
             11'h199: data = 8'b11000110; // **   **
             11'h19a: data = 8'b11000110; // **   **
             11'h19b: data = 8'b01111100; //  *****
             11'h19c: data = 8'b00000000; // 
             11'h19d: data = 8'b00000000; // 
             11'h19e: data = 8'b00000000; // 
             11'h19f: data = 8'b00000000; // 
    
    //code x1a  
             11'h1a0: data = 8'b00000000; // 
             11'h1a1: data = 8'b00000000; // 
             11'h1a2: data = 8'b00111111; // ******
             11'h1a3: data = 8'b01100110; //  **  **
             11'h1a4: data = 8'b01100110; //  **  **
             11'h1a5: data = 8'b01100110; //  **  **
             11'h1a6: data = 8'b01111100; //  *****
             11'h1a7: data = 8'b00001100; //  **
             11'h1a8: data = 8'b00001100; //  **
             11'h1a9: data = 8'b00001100; //  **
             11'h1aa: data = 8'b00001100; //  **
             11'h1ab: data = 8'b00011111; // ****
             11'h1ac: data = 8'b00000000; // 
             11'h1ad: data = 8'b00000000; // 
             11'h1ae: data = 8'b00000000; // 
             11'h1af: data = 8'b00000000; // 
    
    //code x1b
             11'h1b0: data = 8'b00000000; // 
             11'h1b1: data = 8'b00000000; // 
             11'h1b2: data = 8'b01111100; //  *****
             11'h1b3: data = 8'b11000110; // **   **
             11'h1b4: data = 8'b11000110; // **   **
             11'h1b5: data = 8'b11000110; // **   **
             11'h1b6: data = 8'b11000110; // **   **
             11'h1b7: data = 8'b11000110; // **   **
             11'h1b8: data = 8'b11000110; // **   **
             11'h1b9: data = 8'b11010110; // ** * **
             11'h1ba: data = 8'b11011110; // ** ****
             11'h1bb: data = 8'b01111100; //  *****
             11'h1bc: data = 8'b00001100; //     **
             11'h1bd: data = 8'b00001110; //     ***
             11'h1be: data = 8'b00000000; // 
             11'h1bf: data = 8'b00000000; // 
    
    //code x1c   
             11'h1c0: data = 8'b00000000; // 
             11'h1c1: data = 8'b00000000; // 
             11'h1c2: data = 8'b00111111; // ******
             11'h1c3: data = 8'b01100110; //  **  **
             11'h1c4: data = 8'b01100110; //  **  **
             11'h1c5: data = 8'b01100110; //  **  **
             11'h1c6: data = 8'b00111110; //  *****
             11'h1c7: data = 8'b00110110; //  ** **
             11'h1c8: data = 8'b01100110; //  **  **
             11'h1c9: data = 8'b01100110; //  **  **
             11'h1ca: data = 8'b01100110; //  **  **
             11'h1cb: data = 8'b01100111; // ***  **
             11'h1cc: data = 8'b00000000; // 
             11'h1cd: data = 8'b00000000; // 
             11'h1ce: data = 8'b00000000; // 
             11'h1cf: data = 8'b00000000; // 
    
    //code x1d   
             11'h1d0: data = 8'b00000000; // 
             11'h1d1: data = 8'b00000000; // 
             11'h1d2: data = 8'b01111100; //  *****
             11'h1d3: data = 8'b01100011; // **   **
             11'h1d4: data = 8'b01100011; // **   **
             11'h1d5: data = 8'b00000110; //  **
             11'h1d6: data = 8'b00011100; //   ***
             11'h1d7: data = 8'b00110000; //     **
             11'h1d8: data = 8'b01100000; //      **
             11'h1d9: data = 8'b01100011; // **   **
             11'h1da: data = 8'b01100011; // **   **
             11'h1db: data = 8'b00111110; //  *****
             11'h1dc: data = 8'b00000000; // 
             11'h1dd: data = 8'b00000000; // 
             11'h1de: data = 8'b00000000; // 
             11'h1df: data = 8'b00000000; // 
    
    //code x1e   
             11'h1e0: data = 8'b00000000; // 
             11'h1e1: data = 8'b00000000; // 
             11'h1e2: data = 8'b11111111; // ********
             11'h1e3: data = 8'b11011011; // ** ** **
             11'h1e4: data = 8'b10011001; // *  **  *
             11'h1e5: data = 8'b00011000; //    **
             11'h1e6: data = 8'b00011000; //    **
             11'h1e7: data = 8'b00011000; //    **
             11'h1e8: data = 8'b00011000; //    **
             11'h1e9: data = 8'b00011000; //    **
             11'h1ea: data = 8'b00011000; //    **
             11'h1eb: data = 8'b00111100; //   ****
             11'h1ec: data = 8'b00000000; // 
             11'h1ed: data = 8'b00000000; // 
             11'h1ee: data = 8'b00000000; // 
             11'h1ef: data = 8'b00000000; // 
    
    //code x1f   
             11'h1f0: data = 8'b00000000; // 
             11'h1f1: data = 8'b00000000; // 
             11'h1f2: data = 8'b11000110; // **   **
             11'h1f3: data = 8'b11000110; // **   **
             11'h1f4: data = 8'b11000110; // **   **
             11'h515: data = 8'b11000110; // **   **
             11'h1f6: data = 8'b11000110; // **   **
             11'h1f7: data = 8'b11000110; // **   **
             11'h1f8: data = 8'b11000110; // **   **
             11'h1f9: data = 8'b11000110; // **   **
             11'h1fa: data = 8'b11000110; // **   **
             11'h1fb: data = 8'b01111100; //  *****
             11'h1fc: data = 8'b00000000; // 
             11'h1fd: data = 8'b00000000; // 
             11'h1fe: data = 8'b00000000; // 
             11'h1ff: data = 8'b00000000; // 
    
    //code x20 
             11'h200: data = 8'b00000000; // 
             11'h201: data = 8'b00000000; // 
             11'h202: data = 8'b11000011; // **    **
             11'h203: data = 8'b11000011; // **    **
             11'h204: data = 8'b11000011; // **    **
             11'h205: data = 8'b11000011; // **    **
             11'h206: data = 8'b11000011; // **    **
             11'h207: data = 8'b11000011; // **    **
             11'h208: data = 8'b11000011; // **    **
             11'h209: data = 8'b01100110; //  **  **
             11'h20a: data = 8'b00111100; //   ****
             11'h20b: data = 8'b00011000; //    **
             11'h20c: data = 8'b00000000; // 
             11'h20d: data = 8'b00000000; // 
             11'h20e: data = 8'b00000000; // 
             11'h20f: data = 8'b00000000; // 
    
    //code x21   
             11'h210: data = 8'b00000000; // 
             11'h211: data = 8'b00000000; // 
             11'h212: data = 8'b11000011; // **    **
             11'h213: data = 8'b11000011; // **    **
             11'h214: data = 8'b11000011; // **    **
             11'h215: data = 8'b11000011; // **    **
             11'h216: data = 8'b11000011; // **    **
             11'h217: data = 8'b11011011; // ** ** **
             11'h218: data = 8'b11011011; // ** ** **
             11'h219: data = 8'b11111111; // ********
             11'h21a: data = 8'b01100110; //  **  **
             11'h21b: data = 8'b01100110; //  **  **
             11'h21c: data = 8'b00000000; // 
             11'h21d: data = 8'b00000000; // 
             11'h21e: data = 8'b00000000; // 
             11'h21f: data = 8'b00000000; // 
    
    //code x22   
             11'h220: data = 8'b00000000; // 
             11'h221: data = 8'b00000000; // 
             11'h222: data = 8'b11000011; // **    **
             11'h223: data = 8'b11000011; // **    **
             11'h224: data = 8'b01100110; //  **  **
             11'h225: data = 8'b00111100; //   ****
             11'h226: data = 8'b00011000; //    **
             11'h227: data = 8'b00011000; //    **
             11'h228: data = 8'b00111100; //   ****
             11'h229: data = 8'b01100110; //  **  **
             11'h22a: data = 8'b11000011; // **    **
             11'h22b: data = 8'b11000011; // **    **
             11'h22c: data = 8'b00000000; // 
             11'h22d: data = 8'b00000000; // 
             11'h22e: data = 8'b00000000; // 
             11'h22f: data = 8'b00000000; // 
    
    //code x23  
             11'h230: data = 8'b00000000; // 
             11'h231: data = 8'b00000000; // 
             11'h232: data = 8'b11000011; // **    **
             11'h233: data = 8'b11000011; // **    **
             11'h234: data = 8'b11000011; // **    **
             11'h235: data = 8'b01100110; //  **  **
             11'h236: data = 8'b00111100; //   ****
             11'h237: data = 8'b00011000; //    **
             11'h238: data = 8'b00011000; //    **
             11'h239: data = 8'b00011000; //    **
             11'h23a: data = 8'b00011000; //    **
             11'h23b: data = 8'b00111100; //   ****
             11'h23c: data = 8'b00000000; // 
             11'h23d: data = 8'b00000000; // 
             11'h23e: data = 8'b00000000; // 
             11'h23f: data = 8'b00000000; // 
    
    //code x24   
             11'h240: data = 8'b00000000; // 
             11'h241: data = 8'b00000000; // 
             11'h242: data = 8'b11111111; // ********
             11'h243: data = 8'b11000011; // **    **
             11'h244: data = 8'b10000110; // *    **
             11'h245: data = 8'b00001100; //     **
             11'h246: data = 8'b00011000; //    **
             11'h247: data = 8'b00110000; //   **
             11'h248: data = 8'b01100000; //  **
             11'h249: data = 8'b11000001; // **     *
             11'h24a: data = 8'b11000011; // **    **
             11'h24b: data = 8'b11111111; // ********
             11'h24c: data = 8'b00000000; // 
             11'h24d: data = 8'b00000000; // 
             11'h24e: data = 8'b00000000; // 
             11'h24f: data = 8'b00000000; //
             
    //code 25
             11'h250: data = 8'b00000000; // 
             11'h251: data = 8'b00000000; // 
             11'h252: data = 8'b01000010; //  *    *
             11'h253: data = 8'b11100111; // ***  ***
             11'h254: data = 8'b01000010; // ***  ***
             11'h255: data = 8'b00000000; //  *    *
             11'h256: data = 8'b00000000; //   
             11'h257: data = 8'b00000000; //   
             11'h258: data = 8'b00111100; //   ****
             11'h259: data = 8'b01000010; //  *    *
             11'h25a: data = 8'b10000001; // *      *
             11'h25b: data = 8'b10000001; // *      *
             11'h25c: data = 8'b00000000; // 
             11'h25d: data = 8'b00000000; // 
             11'h25e: data = 8'b00000000; // 
             11'h25f: data = 8'b00000000; //
             
			 default: data = 8'b00000000;
    endcase
end

endmodule